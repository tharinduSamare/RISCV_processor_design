module mem_controller 
#(
    ADDRESS_WIDTH = 8,
    DATA_WIDTH = 32
)
(
    input logic clk,wrEn,
    input logic [ADDRESS_WIDTH-1:0]address,
    input logic [DATA_WIDTH-1:0]data

);





endmodule : mem_controller