module top #(

)(
    input logic clk, rstN
);




    
endmodule